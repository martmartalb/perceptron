library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;

entity test_Weights is
--   port (
--     clock
--   ) ;
end test_Weights ; 

architecture arch of test_Weights is

component Bias 
    Generic ( 

    };
    Port (

    );
end component;

end architecture ;