library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package bus_pkg is
    type bus_array is array(natural range <>) of signed;
end package;

package body bus_pkg is

end bus_pkg;